magic
tech scmos
timestamp 1731129436
<< nwell >>
rect -57 44 61 57
rect -57 30 60 44
rect -57 -78 63 30
<< polysilicon >>
rect 11 7 16 10
rect -33 5 -31 6
rect -11 5 -9 6
rect 11 3 14 7
rect 11 1 16 3
rect 36 5 38 8
rect -33 -21 -31 -19
rect -11 -21 -9 -19
rect 11 -22 16 -19
rect 36 -21 38 -19
rect 36 -45 38 -43
rect 36 -72 38 -69
rect -10 -113 -8 -112
rect 18 -113 20 -112
rect 48 -113 50 -112
rect -34 -119 -32 -117
rect -34 -126 -32 -124
rect -10 -125 -8 -123
rect 18 -125 20 -123
rect 48 -125 50 -123
rect -10 -143 -8 -141
rect 18 -143 20 -141
rect 48 -143 50 -141
rect -10 -154 -8 -153
rect 18 -154 20 -153
rect 48 -154 50 -153
<< ndiffusion >>
rect -39 -120 -34 -119
rect -35 -124 -34 -120
rect -32 -124 -27 -119
rect -15 -120 -10 -113
rect -11 -123 -10 -120
rect -8 -123 -3 -113
rect 13 -121 18 -113
rect 17 -123 18 -121
rect 20 -123 25 -113
rect 43 -123 48 -113
rect 50 -116 55 -113
rect 50 -120 53 -116
rect 50 -123 55 -120
rect -11 -145 -10 -143
rect -15 -153 -10 -145
rect -8 -144 -3 -143
rect -8 -148 -5 -144
rect 17 -145 18 -143
rect -8 -153 -3 -148
rect 13 -153 18 -145
rect 20 -145 25 -143
rect 47 -145 48 -143
rect 20 -149 23 -145
rect 20 -153 25 -149
rect 43 -153 48 -145
rect 50 -145 55 -143
rect 50 -149 53 -145
rect 50 -153 55 -149
<< pdiffusion >>
rect -38 -2 -33 5
rect -34 -6 -33 -2
rect -38 -19 -33 -6
rect -31 -19 -26 5
rect -16 -2 -11 5
rect -12 -6 -11 -2
rect -16 -19 -11 -6
rect -9 -19 -4 5
rect 35 2 36 5
rect 6 -2 11 1
rect 10 -6 11 -2
rect 6 -19 11 -6
rect 16 0 21 1
rect 16 -4 18 0
rect 16 -19 21 -4
rect 31 -19 36 2
rect 38 -19 43 5
rect 31 -69 36 -45
rect 38 -50 43 -45
rect 38 -54 40 -50
rect 38 -63 43 -54
rect 38 -67 41 -63
rect 38 -69 43 -67
<< metal1 >>
rect -29 6 -11 9
rect 18 0 21 6
rect 40 -25 54 -22
rect 11 -40 16 -26
rect 11 -43 36 -40
rect 51 -51 54 -25
rect 44 -54 54 -51
rect -39 -94 58 -91
rect -34 -113 -31 -94
rect -10 -108 -7 -94
rect 18 -108 21 -94
rect 48 -108 51 -94
rect -10 -165 -7 -158
rect 18 -165 21 -158
rect 48 -165 51 -158
rect -23 -169 63 -165
<< metal2 >>
rect -43 38 60 44
rect -50 35 60 38
rect -50 -2 -44 35
rect -20 -2 -17 35
rect -50 -6 -35 -2
rect -20 -5 -13 -2
rect 2 -3 5 35
rect 31 2 34 35
rect 2 -6 8 -3
rect -28 -41 -25 -17
rect -50 -44 -25 -41
rect -50 -124 -47 -44
rect 41 -67 49 -64
rect 46 -81 49 -67
rect 45 -84 49 -81
rect 37 -87 48 -84
rect 37 -117 40 -87
rect 37 -120 46 -117
rect 53 -120 62 -117
rect -40 -124 -36 -122
rect -50 -125 -36 -124
rect -50 -127 -37 -125
rect -40 -128 -37 -127
rect -15 -145 -11 -120
rect 13 -145 16 -121
rect 59 -130 62 -120
rect 43 -133 62 -130
rect 43 -145 46 -133
rect -5 -148 5 -145
rect 2 -202 5 -148
rect 23 -149 33 -145
rect 53 -147 63 -146
rect 53 -149 64 -147
rect 30 -202 33 -149
rect 60 -200 64 -149
rect 59 -202 64 -200
rect -24 -203 64 -202
rect -24 -206 62 -203
<< ntransistor >>
rect -34 -124 -32 -119
rect -10 -123 -8 -113
rect 18 -123 20 -113
rect 48 -123 50 -113
rect -10 -153 -8 -143
rect 18 -153 20 -143
rect 48 -153 50 -143
<< ptransistor >>
rect -33 -19 -31 5
rect -11 -19 -9 5
rect 11 -19 16 1
rect 36 -19 38 5
rect 36 -69 38 -45
<< polycontact >>
rect -33 6 -29 10
rect -11 6 -7 10
rect 14 3 18 7
rect 11 -26 16 -22
rect 36 -25 40 -21
rect 36 -43 40 -39
rect -10 -112 -6 -108
rect 18 -112 22 -108
rect 48 -112 52 -108
rect -34 -117 -30 -113
rect -10 -158 -6 -154
rect 18 -158 22 -154
rect 48 -158 52 -154
<< ndcontact >>
rect -39 -124 -35 -120
rect -15 -124 -11 -120
rect 13 -125 17 -121
rect 53 -120 57 -116
rect -15 -145 -11 -141
rect -5 -148 -1 -144
rect 13 -145 17 -141
rect 43 -145 47 -141
rect 23 -149 27 -145
rect 53 -149 57 -145
<< pdcontact >>
rect -38 -6 -34 -2
rect -16 -6 -12 -2
rect 31 2 35 6
rect 6 -6 10 -2
rect 18 -4 22 0
rect 40 -54 44 -50
rect 41 -67 45 -63
<< end >>
